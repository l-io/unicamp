* C:\Users\Squadra\Desktop\ee610\sim2\sim2.sch

* Schematics Version 9.1 - Web Update 1
* Fri Jan 22 15:28:45 2021



** Analysis setup **
.tran 0ns 1000ns 970ns 0.1ps
.OP 
.LIB "C:\Users\Squadra\Desktop\ee610\sim1\sim1.lib"


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "sim2.net"
.INC "sim2.als"


.probe


.END
